*** SPICE deck for cell osc11{sch} from library lab1
*** Created on Wed Feb 05, 2020 22:48:40
*** Last revised on Wed Feb 05, 2020 22:54:18
*** Written on Wed Feb 05, 2020 23:26:26 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include C:\Users\12217\Documents\GitHub\1920SemB_EE4204_RayC\lab1\scmos18.txt

*** SUBCIRCUIT lab1__inv FROM CELL inv{sch}
.SUBCKT lab1__inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.2U W=0.9U
Mpmos@1 vdd in out vdd P L=0.2U W=1.8U
.ENDS lab1__inv

.global gnd vdd ring_out_11

*** TOP LEVEL CELL: osc11{sch}
Xinv@0 ring_out_11 net@0 lab1__inv
Xinv@1 net@0 net@11 lab1__inv
Xinv@2 net@11 net@2 lab1__inv
Xinv@3 net@2 net@3 lab1__inv
Xinv@4 net@3 net@27 lab1__inv
Xinv@5 net@26 net@15 lab1__inv
Xinv@6 net@15 net@17 lab1__inv
Xinv@7 net@17 net@19 lab1__inv
Xinv@8 net@19 net@22 lab1__inv
Xinv@9 net@22 ring_out_11 lab1__inv
Xinv@10 net@27 net@26 lab1__inv
* Trailer cards are described in this file:
.include C:\Users\12217\Documents\GitHub\1920SemB_EE4204_RayC\lab1\user_append.spi
.END
